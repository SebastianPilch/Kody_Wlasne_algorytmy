`timescale 1ns / 1ps
//-----------------------------------------------
// Company: agh
//-----------------------------------------------
module i_mem
(
  input [7:0]address,
  output [31:0]data
);
//-----------------------------------------------
//instruction memory
wire [31:0]program[255:0];
reg Rx = 4'h1;
reg Rd = 4'h2;

////


//////////////////////////////////////////////////
//  |___  |  / ___ \  |  _ \      /     |
//     / /  | |   | | | | \ |    /__/|  |
//    / /   | |___| | | |  ||        |  |
//   / /__  |  ___  | | |_/ |       _|  |_
//  |_____| |_|   |_| |____/       |______|
////////////////////////////////////////////////////////
//TESTY MOV i MOVI
// zadanie 13.1
// na zmian� wpisuje warto�ci 2 i 4 do R1
// nast�pnie przepisuje warto�� z R1 do R2 
// a nast�pnie si� zap�tla poprzez jumpi
///




//assign program[0] = 32'b00000000000101101000000100000100; //movi R1, 4, 
//assign program[1] = 32'b00000000000100010110001000000000; // //mov R1, R2, 
//assign program[2] = 32'b00000000000101101000000100000010; //movi R1, 2, 
//assign program[3] = 32'b00000000000100010110001000000000; // //movi R1, R2, 
//assign program[4] = 32'b00000001001100101000001100000000; //jumpi 0


//////////////////////////////////////////////////
//  |___  |  / ___ \  |  _ \      /   _   \
//     / /  | |   | | | | \ |    |__/ /  /
//    / /   | |___| | | |  ||        /  /
//   / /__  |  ___  | | |_/ |       /  /___
//  |_____| |_|   |_| |____/       |_______|
////////////////////////////////////////////////////////
////
//TESTY add, addi inwencja tw�rcza moja do usuni�cia 
// testy add i addi przy okazji nop i jnz
// stworzenie p�tli czekaj�cej 5ns*16
// wykonanie inkrementacja R2 poprzez addi
///
//assign program[0] = 32'b00000000000101101000000000000011;//movi R0, 0x03 
//assign program[1] = 32'b00000000000101101000000100010000;//movi R1, 0x10
//assign program[2] = 32'b00000000000100000001001000000000;//add R2, R0, R1
//assign program[3] = 32'b00000000000100001000001100100000;//addi R3, R0, 0x20
//assign program[4] = 32'b00000000000101101000010011101111;//movi R4, 0xef
//assign program[5] = 32'b00000000000101100000000000000000;//nop 
//assign program[6] = 32'b00000000000101100000000000000000;//nop 
//assign program[7] = 32'b00000000000101100000000000000000;//nop 
//assign program[8] = 32'b00000000000101001000010000000001;//addi R4, R4, 0x01
//assign program[9] = 32'b00000011001101001110011100000101;//jnz R4, 0x05



//////////////////////////////////////////////////
//  |___  |  / ___ \  |  _ \      /   _   \
//     / /  | |   | | | | \ |    |__/ /  /
//    / /   | |___| | | |  ||      __ \  \
//   / /__  |  ___  | | |_/ |    /  /_/   |
//  |_____| |_|   |_| |____/     \_______/
////////////////////////////////////////////////////////
////
//ZADANIE 13.5
//  Tre�� w zadaniu na upelu
///

assign program[0] = 32'b00000000000101101000000000000000;//movi R0, 0x00
assign program[1] = 32'b00000000000101101000000100000100;//movi R1, 0x04
assign program[2] = 32'b00000000000100001000000000000001;//addi R0, R0, 0x01
assign program[3] = 32'b00000000000000000001101000000000;//and R2, R0, R1
assign program[4] = 32'b00000010001100101110011100000010;//jz R2, 0x02
assign program[5] = 32'b00000000000101101000001100000001;//movi R3, 0x01


//////////////////////////////////////////////////
//  |___  |  / ___ \  |  _ \      /   _  |
//     / /  | |   | | | | \ |    |  /__| |
//    / /   | |___| | | |  ||    |____   |
//   / /__  |  ___  | | |_/ |         |  |
//  |_____| |_|   |_| |____/          |__| 
////////////////////////////////////////////////////////
////
//ZADANIE 14.1
//  Tre�� w zadaniu na upelu
///


//assign program[0] = 32'b00000000000101101000100000000000;//loadi R0, 0x00  #0
//assign program[1] = 32'b00000000000101101000100100000001;//loadi R1, 0x01   #1 
//assign program[2] = 32'b00000000000101101000101000000010;//loadi R2, 0x02  #2
//assign program[3] = 32'b00000000000101101000001100000110;//movi R3, 0x06   #3
//assign program[4] = 32'b00000000000101101000010100000001;//movi R5, 0x01   #4
//assign program[5] = 32'b00000001000101101110011100010000;//jumpi 0x10 1s  #5
//assign program[6] = 32'b00000000000101101000010100000010;//movi R5, 0x02   #6
//assign program[7] = 32'b00000000000001001000001100000001;//andi R3, R4, 0x01  #7
//assign program[8] = 32'b00000011001100111110011100000111;//jnz R3, 0x07  #8
//assign program[9] = 32'b00000000000101101000001100001100;//movi R3, 0x0c   #9
//assign program[10] = 32'b00000000000101101000010100000100;//movi R5, 0x04  #10
//assign program[11] = 32'b00000001000101101110011100010000;//jumpi 0x10 1s  #11
//assign program[12] = 32'b00000000000101101000010100001000;//movi R5, 0x08  #12
//assign program[13] = 32'b00000000000001001000001100000010;//andi R3, R4, 0x10  #13
//assign program[14] = 32'b00000011001100111110011100001101;//jnz R3, 0x0d  #14
//assign program[15] = 32'b00000001000101101110011100000011;//jumpi 0x03  #15
//assign program[16] = 32'b00000000000100001000000000000001;//addi R0, R0, 0x01   #16
//assign program[17] = 32'b00000011001100001110011100010000;//jnz R0, 0x10        #17
//assign program[18] = 32'b00000000000101101000100000000000;//loadi R0, 0x00      #18
//assign program[19] = 32'b00000000000100011000000100000001;//addi R1, R1, 0x01   #19
//assign program[20] = 32'b00000000000101100000000000000000;//nop    		    #20
//assign program[21] = 32'b00000011001100011110011100010000;//jnz R1, 0x10        #21
//assign program[22] = 32'b00000000000101101000100100000001;//loadi R1, 0x01      #22
//assign program[23] = 32'b00000000000100101000001000000001;//addi R2, R2, 0x01   #23
//assign program[24] = 32'b00000000000101100000000000000000;//nop    	 	    #24
//assign program[25] = 32'b00000011001100101110011100010000;//jnz R2, 0x10   	    #25
//assign program[26] = 32'b00000000000101101000101000000010;//loadi R2, 0x02      #26
//assign program[27] = 32'b00000001000101100011011100000000;//jump R3   	    #27

//////////////////////////////////////////////////
//  |___  |  / ___ \  |  _ \      |   ___|
//     / /  | |   | | | | \ |     |  /___
//    / /   | |___| | | |  ||     \____  \
//   / /__  |  ___  | | |_/ |      ____\  |
//  |_____| |_|   |_| |____/      |______/      
////////////////////////////////////////////////////////
////
//ZADANIE 14.1
//  �le zrobione 14.1 ale mo�e wyjdzie fajnie
///

//assign program[0] = 32'b00000000000101101000010100000011;//movi R5, 0x03 
//assign program[1] = 32'b00000000000101101000100000000000;//loadi R0, 0x00
//assign program[2] = 32'b00000000000101101000100100000001;//loadi R1, 0x01
//assign program[3] = 32'b00000000000101101000101000000010;//loadi R2, 0x02
//assign program[4] = 32'b00000000000100001000000000000001;//addi R0, R0, 0x01
//assign program[5] = 32'b00000011001100001110011100000100;//jnz R0, 0x04
//assign program[6] = 32'b00000000000101101000100000000000;//loadi R0, 0x00
//assign program[7] = 32'b00000000000100011000000100000001;//addi R1, R1, 0x01
//assign program[8] = 32'b00000000000101100000000000000000;//nop 
//assign program[9] = 32'b00000011001100011110011100000100;//jnz R1, 0x04
//assign program[10] = 32'b00000000000101101000100100000001;//loadi R1, 0x01
//assign program[11] = 32'b00000000000100101000001000000001;//addi R2, R2, 0x01
//assign program[12] = 32'b00000000000101100000000000000000;//nop 
//assign program[13] = 32'b00000011001100101110011100000100;//jnz R2, 0x04
//assign program[14] = 32'b00000000000101100000000000000000;//nop 
//assign program[15] = 32'b00000000000101100000000000000000;//nop 
//assign program[16] = 32'b00000000000101101000101000000010;//loadi R2, 0x02 
//assign program[17] = 32'b00000000000101010101010100000000;//add R5, R5, R5
//assign program[18] = 32'b00000000000100001000000000000001;//addi R0, R0, 0x01
//assign program[19] = 32'b00000011001100001110011100010011;//jnz R0, 0x13
//assign program[20] = 32'b00000000000101101000100000000000;//loadi R0, 0x00
//assign program[21] = 32'b00000000000100011000000100000001;//addi R1, R1, 0x01
//assign program[22] = 32'b00000000000101100000000000000000;//nop 
//assign program[23] = 32'b00000011001100011110011100000100;//jnz R1, 0x04
//assign program[24] = 32'b00000000000101101000100100000001;//loadi R1, 0x01
//assign program[25] = 32'b00000000000100101000001000000001;//addi R2, R2, 0x01
//assign program[26] = 32'b00000000000101100000000000000000;//nop 
//assign program[27] = 32'b00000011001100101110011100010011;//jnz R2, 0x13
//assign program[28] = 32'b00000000000101101000101000000010;//loadi R2, 0x02 
//assign program[29] = 32'b00000000000101000100010000000000;//add R4, R4, R4 
//assign program[30] = 32'b00000000000101011000010100000001;//addi R5, R5, 0x01
//assign program[31] = 32'b00000001000101101110011100010011;//jumpi 0x13



//-----------------------------------------------
assign data=program[address];
//-----------------------------------------------
endmodule
//-----------------------------------------------